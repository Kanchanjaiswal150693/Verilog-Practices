module ModuleDwithDelay_tb;
  reg a,b,c;
  wire out;
  
  ModuleDwithDelay DelayD(out,a,b,c);
  initial
  begin
    a=1'b0;
    b=1'b0;
    c=1'b0;
    #10;
    a=1'b1;
    b=1'b1;
    c=1'b1;
    #10;
    a=1'b1;
    b=1'b0;
    c=1'b0;
    
  end
endmodule 
