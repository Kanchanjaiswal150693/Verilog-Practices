module mynor(out,a,b);
  output out;
  input a,b;
  
  nor nor1(out,a,b);
  
endmodule
