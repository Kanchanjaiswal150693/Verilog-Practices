module my_invertor(y,a);
  input a;
  output y;
  //initial begin
    assign y=~a;
  //end
  
endmodule

  
