module myxor(out,a,b);
  output out;
  input a,b;
  
  xor myxor1(out,a,b);
  
endmodule
