module my_and(out, a, b);
  output out;
  input a, b;
  
  and and1(out, a, b);
  
endmodule
