module myxnor(out,a,b);
  output out;
  input a,b;
  
  xnor myxnor1(out,a,b);
  
endmodule
