module my_or(out,a,b);
  output out;
  input a,b;
  
  or myor1(out,a,b);
  
endmodule
