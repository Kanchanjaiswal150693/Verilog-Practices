module TwoinOneMultiplexerusingDFM()
